module LSU
(
input [31:0] addr,
input [31:0] wdata,

output [23:0] addr_1,
output [23:0] addr_2,

output [31:0] out_1,
output [31:0] out_2
);

generate

endgenerate

endmodule