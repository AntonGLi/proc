module core (
input logic         clk_i,
input logic         rst_i,
input logic  [31:0] instr_i,
input logic  [31:0] mem_rd_i,
output logic        mem_wd_o,
output logic        mem_we_o,
output logic        mem_addr_o,
output logic [2:0]  mem_size_o,
output logic        mem_req_o,
output logic [31:0] instr_addr_o,
);

//instruction address (pc)
logic [31:0] pc;
logic [31:0] pc_next;
logic pc_en;

always_ff @(posedge clk) begin
  if (rst) begin
    pc = '0;
  end else begin
    if (pc_en) begin
      pc = pc_next;
    end
  end
end

assign instr_addr_o = pc;

//decoding instruction
logic [31:0] fetched_instr;

assign fetched_instr = instr_i;

  //defining constants
logic [11:0] cI, [31:0] I;
logic [11:0] cS, [31:0] S;
logic [12:0] cB, [31:0] B;
logic [20:0] cJ, [31:0] J;
logic [19:0] cU, [31:0] U;

  //from instr
assign cI =   fetched_instr[31:20];
assign cS = {
              fetched_instr[31:25], 
              fetched_instr[11:7]
            };
assign cB = {
              fetched_instr[31], 
              fetched_instr[7], 
              fetched_instr[30:25], 
              fetched_instr[11:8], 
              1'b0
            };
assign cJ = {
              fetched_instr[31], 
              fetched_instr[19:12], 
              fetched_instr[20], 
              fetched_instr[30:21], 
              1'b0
            };
assign cU =   fetched_instr[31:12];

  //to 32 bit
assign  I = {20{cI[11]}, cI};
assign  S = {20{cS[11]}, cS};
assign  B = {19{cB[12]}, cB};
assign  J = {11{cJ[20]}, cJ};
assign  U = {cU, 12'b0};

//control signals
logic [1:0]   a_sel;
logic [2:0]   b_sel;
logic [4:0]   alu_op;
logic [2:0]   csr_op;
logic         csr_we;
logic         mem_req;
logic         mem_we;
logic [2:0]   mem_size;
logic         gpr_we;
logic [1:0]   wb_sel;
logic         illegal_instr;
logic         branch;
logic         jal;
logic         jalr;
logic         mret;

assign mem_we_o   = mem_we;
assign mem_size_o = mem_size;
assign mem_req_o  = mem_req;
assign pc_en = illegal_instr;

//decoder
decoder dc1 (
.fetched_instr_i  (fetched_instr),
.a_sel_o          (a_sel),
.b_sel_o          (b_sel),
.alu_op_o         (oper),
.csr_op_o         (csr_oper),
.csr_we_o         (csr_we),
.mem_req_o        (mem_req),
.mem_we_o         (mem_we),
.mem_size_o       (mem_size),
.gpr_we_o         (gpr_we),
.wb_sel_o         (wb_sel),
.illegal_instr_o  (illegal_instr),
.branch_o         (branch),
.jal_o            (jal),
.jalr_o           (jalr),
.mret_o           (mret)
);

//reg file ports and connect
logic [4:0]   ra1; 
logic [4:0]   ra2; 
logic [4:0]   wa; 
logic         we; 
logic [31:0]  wdata; 
logic [31:0]  rd1; 
logic [31:0]  rd2;

always_comb begin
  we  = gpr_we;
  ra1 = fetched_instr[19:15];
  ra2 = fetched_instr[24:20];
  wa  = fetched_instr[11:7];
  case (wb_sel)
    2'd0: wdata = alu_res;
    2'd1: wdata = mem_rd_i;
    default: wdata = '0;
  endcase
end

Register_file meme1 (
  .clk(clk),

  .WrEn(we),
  .upr_in(wa),
  .in(wdata),

  .upr_A(ra1),
  .upr_B(ra2),

  .A(rd1),
  .B(rd2)
);

//alu
logic [31:0] alu_a;
logic [31:0] alu_b;
logic [4:0]  alu_oper;
logic [31:0] alu_res, 
logic flag;

always_comb begin
  oper = alu_op;
  case (a_sel)
    2'd0:     a = rd1;
    2'd1:     a = pc;
    2'd2:     a = '0;
    default:  a = '0;
  endcase
  case (b_sel)
    3'd0:     b = rd2;
    3'd1:     b = I;
    3'd2:     b = U;
    3'd3:     b = S;
    3'd4:     b = 32'd4;
  endcase
end

ALU alu1 (
  .A(alu_a),
  .B(alu_b),
  .Upr_ALU(alu_oper),
  .C(flag),
  .Out_ALU(alu_res)
);

//pc logic
logic [31:0] I_addr;
logic [31:0] bj;
logic [31:0] bj4;
logic [31:0] bj4_addr;
logic        bj_sel;
logic        bj4_sel;

assign I_addr = rd1 + I;
assign bj4_addr = bj4 + pc;

assign bj_sel   = b;
assign bj4_sel  = jal | (flag & b);

mux2 mux_bj (
.a_1(B),
.b_0(J),
.sel(bj_sel),
.c(bj)
);

mux2 mux_bj4 (
.a_1(bj),
.b_0(32'd4),
.sel(bj4_sel),
.c(bj4)
);

mux2 mux_pc_next (
.a_1(I_addr),
.b_0(bj4_addr),
.sel(jalr),
.c(pc_next)
);

endmodule

